`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company:
// Engineer:
//
// Create Date:
// Design Name:
// Module Name: ShiftLogical
// Project Name:
// Target Devices:
// Tool Versions:
// Description:
//
// Dependencies:
//
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
//
//////////////////////////////////////////////////////////////////////////////////


module ShiftLogical (
    input  [31:0] in1,  //输入1
    input  [31:0] in2,  //输入2
    input  [ 1:0] sel,  //运算选择
    output [31:0] out   //运算结果
);

endmodule
